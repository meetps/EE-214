library verilog;
use verilog.vl_types.all;
entity sram is
end sram;
